module(ouput y, input a);
  assign y= ~a;
endmodule
